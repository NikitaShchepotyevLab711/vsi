module xci2_buf (
    input wire a,
    output wire y
);

assign y = a;    

endmodule